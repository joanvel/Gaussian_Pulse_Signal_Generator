library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity LUT is
	generic(g_bits:integer:=16
				;g_lines:integer:=11);
	port
			(i_Data:in std_logic_vector(g_lines-1 downto 0)
			;o_Data:out std_logic_vector(g_bits-1 downto 0)
			);
end LUT;

Architecture RTL of LUT is
	type exp is array (0 to 2**(g_lines)-1) of integer;
	constant values: exp:=(1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3
									,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4
									,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7
									,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,11
									,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14
									,14,14,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,17,17,17,17,17,17,17,18,18,18,18,18,18,19,19,19
									,19,19,19,19,20,20,20,20,20,20,21,21,21,21,21,22,22,22,22,22,22,23,23,23,23,23,24,24,24,24,24,25,25
									,25,25,25,26,26,26,26,27,27,27,27,27,28,28,28,28,29,29,29,29,30,30,30,30,31,31,31,31,32,32,32,32,33
									,33,33,33,34,34,34,34,35,35,35,36,36,36,36,37,37,37,38,38,38,39,39,39,40,40,40,40,41,41,41,42,42,42
									,43,43,43,44,44,45,45,45,46,46,46,47,47,47,48,48,49,49,49,50,50,51,51,51,52,52,53,53,53,54,54,55,55
									,55,56,56,57,57,58,58,59,59,59,60,60,61,61,62,62,63,63,64,64,65,65,66,66,67,67,68,68,69,69,70,70,71
									,71,72,73,73,74,74,75,75,76,76,77,78,78,79,79,80,81,81,82,82,83,84,84,85,86,86,87,88,88,89,89,90,91
									,92,92,93,94,94,95,96,96,97,98,99,99,100,101,101,102,103,104,105,105,106,107,108,108,109,110,111,112
									,112,113,114,115,116,117,117,118,119,120,121,122,123,124,124,125,126,127,128,129,130,131,132,133,134
									,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,159,160
									,161,162,163,164,165,167,168,169,170,171,173,174,175,176,177,179,180,181,182,184,185,186,188,189,190
									,192,193,194,196,197,198,200,201,202,204,205,207,208,209,211,212,214,215,217,218,220,221,223,224,226
									,227,229,230,232,234,235,237,238,240,242,243,245,247,248,250,252,253,255,257,258,260,262,264,266,267
									,269,271,273,275,276,278,280,282,284,286,288,290,291,293,295,297,299,301,303,305,307,309,311,313,315
									,318,320,322,324,326,328,330,332,335,337,339,341,343,346,348,350,353,355,357,359,362,364,367,369,371
									,374,376,379,381,383,386,388,391,393,396,398,401,404,406,409,411,414,417,419,422,425,427,430,433,436
									,438,441,444,447,450,452,455,458,461,464,467,470,473,476,479,482,485,488,491,494,497,500,503,506,510
									,513,516,519,522,526,529,532,536,539,542,546,549,552,556,559,563,566,570,573,577,580,584,587,591,595
									,598,602,605,609,613,617,620,624,628,632,636,639,643,647,651,655,659,663,667,671,675,679,683,687,691
									,696,700,704,708,712,717,721,725,730,734,738,743,747,752,756,761,765,770,774,779,783,788,793,797,802
									,807,811,816,821,826,831,835,840,845,850,855,860,865,870,875,880,885,891,896,901,906,911,917,922,927
									,933,938,943,949,954,960,965,971,976,982,988,993,999,1005,1010,1016,1022,1028,1033,1039,1045,1051
									,1057,1063,1069,1075,1081,1087,1093,1100,1106,1112,1118,1125,1131,1137,1144,1150,1156,1163,1169,1176
									,1182,1189,1196,1202,1209,1216,1222,1229,1236,1243,1250,1256,1263,1270,1277,1284,1291,1299,1306,1313
									,1320,1327,1334,1342,1349,1356,1364,1371,1379,1386,1394,1401,1409,1417,1424,1432,1440,1447,1455,1463
									,1471,1479,1487,1495,1503,1511,1519,1527,1535,1543,1552,1560,1568,1577,1585,1593,1602,1610,1619,1627
									,1636,1645,1653,1662,1671,1680,1688,1697,1706,1715,1724,1733,1742,1751,1761,1770,1779,1788,1798,1807
									,1816,1826,1835,1845,1854,1864,1874,1883,1893,1903,1912,1922,1932,1942,1952,1962,1972,1982,1992,2003
									,2013,2023,2033,2044,2054,2064,2075,2085,2096,2107,2117,2128,2139,2149,2160,2171,2182,2193,2204,2215
									,2226,2237,2249,2260,2271,2282,2294,2305,2317,2328,2340,2351,2363,2375,2386,2398,2410,2422,2434,2446
									,2458,2470,2482,2494,2506,2519,2531,2543,2556,2568,2581,2593,2606,2618,2631,2644,2657,2670,2682,2695
									,2708,2721,2735,2748,2761,2774,2787,2801,2814,2828,2841,2855,2868,2882,2896,2909,2923,2937,2951,2965
									,2979,2993,3007,3021,3036,3050,3064,3079,3093,3108,3122,3137,3151,3166,3181,3196,3211,3226,3241,3256
									,3271,3286,3301,3316,3332,3347,3362,3378,3393,3409,3425,3440,3456,3472,3488,3504,3520,3536,3552,3568
									,3584,3600,3617,3633,3650,3666,3683,3699,3716,3733,3749,3766,3783,3800,3817,3834,3851,3869,3886,3903
									,3920,3938,3955,3973,3991,4008,4026,4044,4062,4079,4097,4115,4134,4152,4170,4188,4206,4225,4243,4262
									,4280,4299,4318,4336,4355,4374,4393,4412,4431,4450,4469,4489,4508,4527,4547,4566,4586,4605,4625,4645
									,4665,4684,4704,4724,4744,4765,4785,4805,4825,4846,4866,4887,4907,4928,4948,4969,4990,5011,5032,5053
									,5074,5095,5116,5138,5159,5180,5202,5223,5245,5266,5288,5310,5332,5354,5376,5398,5420,5442,5464,5487
									,5509,5531,5554,5576,5599,5622,5645,5667,5690,5713,5736,5759,5782,5806,5829,5852,5876,5899,5923,5946
									,5970,5994,6018,6042,6066,6090,6114,6138,6162,6186,6211,6235,6260,6284,6309,6334,6358,6383,6408,6433
									,6458,6483,6508,6533,6559,6584,6610,6635,6661,6686,6712,6738,6764,6790,6815,6842,6868,6894,6920,6946
									,6973,6999,7026,7052,7079,7106,7132,7159,7186,7213,7240,7267,7295,7322,7349,7377,7404,7432,7459,7487
									,7515,7542,7570,7598,7626,7654,7682,7711,7739,7767,7796,7824,7853,7881,7910,7939,7968,7996,8025,8054
									,8083,8113,8142,8171,8201,8230,8259,8289,8319,8348,8378,8408,8438,8468,8498,8528,8558,8588,8619,8649
									,8679,8710,8740,8771,8802,8833,8863,8894,8925,8956,8987,9018,9050,9081,9112,9144,9175,9207,9238,9270
									,9302,9334,9366,9398,9430,9462,9494,9526,9558,9591,9623,9655,9688,9721,9753,9786,9819,9852,9885,9918
									,9951,9984,10017,10050,10083,10117,10150,10184,10217,10251,10285,10318,10352,10386,10420,10454,10488
									,10522,10556,10591,10625,10659,10694,10728,10763,10797,10832,10867,10901,10936,10971,11006,11041
									,11076,11112,11147,11182,11217,11253,11288,11324,11359,11395,11431,11466,11502,11538,11574,11610
									,11646,11682,11718,11754,11791,11827,11863,11900,11936,11973,12010,12046,12083,12120,12157,12193
									,12230,12267,12304,12342,12379,12416,12453,12491,12528,12565,12603,12640,12678,12716,12753,12791
									,12829,12867,12905,12943,12981,13019,13057,13095,13133,13171,13210,13248,13287,13325,13364,13402
									,13441,13479,13518,13557,13596,13634,13673,13712,13751,13790,13829,13869,13908,13947,13986,14026
									,14065,14104,14144,14183,14223,14262,14302,14342,14381,14421,14461,14501,14541,14581,14621,14661
									,14701,14741,14781,14821,14861,14902,14942,14982,15023,15063,15104,15144,15185,15225,15266,15306
									,15347,15388,15429,15469,15510,15551,15592,15633,15674,15715,15756,15797,15838,15879,15920,15962
									,16003,16044,16085,16127,16168,16209,16251,16292,16334,16375,16417,16458,16500,16542,16583,16625
									,16667,16709,16750,16792,16834,16876,16918,16960,17001,17043,17085,17127,17169,17211,17254,17296
									,17338,17380,17422,17464,17506,17549,17591,17633,17675,17718,17760,17802,17845,17887,17929,17972
									,18014,18057,18099,18142,18184,18227,18269,18312,18354,18397,18439,18482,18524,18567,18610,18652
									,18695,18738,18780,18823,18866,18908,18951,18994,19036,19079,19122,19165,19207,19250,19293,19336
									,19378,19421,19464,19507,19549,19592,19635,19678,19721,19763,19806,19849,19892,19935,19977,20020
									,20063,20106,20149,20191,20234,20277,20320,20362,20405,20448,20491,20533,20576,20619,20662,20704
									,20747,20790,20832,20875,20918,20961,21003,21046,21088,21131,21174,21216,21259,21301,21344,21387
									,21429,21472,21514,21557,21599,21642,21684,21726,21769,21811,21854,21896,21938,21980,22023,22065
									,22107,22149,22192,22234,22276,22318,22360,22402,22444,22486,22528,22570,22612,22654,22696,22738
									,22780,22822,22863,22905,22947,22989,23030,23072,23113,23155,23197,23238,23280,23321,23362,23404
									,23445,23486,23528,23569,23610,23651,23692,23733,23774,23815,23856,23897,23938,23979,24020,24060
									,24101,24142,24182,24223,24263,24304,24344,24385,24425,24465,24506,24546,24586,24626,24666,24706
									,24746,24786,24826,24866,24905,24945,24985,25024,25064,25103,25143,25182,25221,25261,25300,25339
									,25378,25417,25456,25495,25534,25573,25611,25650,25689,25727,25766,25804,25843,25881,25919,25957
									,25995,26033,26071,26109,26147,26185,26223,26260,26298,26336,26373,26410,26448,26485,26522,26559
									,26596,26633,26670,26707,26744,26780,26817,26853,26890,26926,26962,26999,27035,27071,27107,27143
									,27179,27214,27250,27286,27321,27357,27392,27427,27462,27497,27532,27567,27602,27637,27672,27706
									,27741,27775,27810,27844,27878,27912,27946,27980,28014,28048,28081,28115,28148,28182,28215,28248
									,28281,28314,28347,28380,28412,28445,28478,28510,28542,28575,28607,28639,28671,28703,28734,28766
									,28798,28829,28860,28892,28923,28954,28985,29016,29046,29077,29108,29138,29168,29199,29229,29259
									,29289,29319,29348,29378,29407,29437,29466,29495,29524,29553,29582,29611,29640,29668,29697,29725
									,29753,29781,29809,29837,29865,29892,29920,29947,29975,30002,30029,30056,30083,30109,30136,30162
									,30189,30215,30241,30267,30293,30319,30345,30370,30396,30421,30446,30471,30496,30521,30546,30570
									,30595,30619,30643,30667,30691,30715,30739,30762,30786,30809,30832,30856,30879,30901,30924,30947
									,30969,30991,31014,31036,31058,31080,31101,31123,31144,31166,31187,31208,31229,31249,31270,31291
									,31311,31331,31351,31371,31391,31411,31431,31450,31469,31489,31508,31527,31545,31564,31582,31601
									,31619,31637,31655,31673,31691,31708,31726,31743,31760,31777,31794,31811,31827,31844,31860,31876
									,31892,31908,31924,31940,31955,31970,31986,32001,32016,32030,32045,32060,32074,32088,32102,32116
									,32130,32143,32157,32170,32184,32197,32209,32222,32235,32247,32260,32272,32284,32296,32308,32319
									,32331,32342,32353,32364,32375,32386,32396,32407,32417,32427,32437,32447,32457,32466,32476,32485
									,32494,32503,32512,32521,32529,32538,32546,32554,32562,32570,32577,32585,32592,32599,32606,32613
									,32620,32626,32633,32639,32645,32651,32657,32663,32668,32674,32679,32684,32689,32694,32698,32703
									,32707,32711,32715,32719,32723,32726,32730,32733,32736,32739,32742,32745,32747,32749,32752,32754
									,32756,32757,32759,32760,32762,32763,32764,32765,32765,32766,32766,32766,32767);
begin
	o_Data <= std_logic_vector(to_unsigned(values(to_integer(unsigned(i_Data))),g_bits));
end RTL;