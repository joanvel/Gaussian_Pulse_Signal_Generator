library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity LUT is
	generic(g_bits:integer:=16
				;g_lines:integer:=8);
	port
			(i_Data:in std_logic_vector(g_lines-1 downto 0)
			;o_Data:out std_logic_vector(g_bits-1 downto 0)
			);
end LUT;

Architecture RTL of LUT is
	type exp is array (0 to 2**(g_lines)-1) of integer;
	constant values: exp:=(0,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,3,3,3,3,
									4,4,4,4,5,5,6,6,7,7,8,8,9,9,10,11,12,12,
									13,14,15,16,17,18,20,21,22,24,26,27,29,
									31,33,35,37,39,42,45,47,50,53,57,60,64,
									67,71,76,80,85,90,95,100,106,112,118,125,
									132,139,147,155,163,172,181,191,201,212,
									223,234,246,259,272,286,301,316,332,348,
									365,383,402,421,441,462,484,507,530,555,
									580,607,635,663,693,724,756,789,823,859,
									895,934,973,1014,1056,1100,1145,1191,1239,
									1289,1340,1393,1448,1504,1562,1621,1683,
									1746,1811,1878,1947,2017,2090,2164,2241,
									2319,2400,2483,2567,2654,2743,2834,2927,
									3023,3120,3220,3322,3426,3532,3640,3751,
									3864,3979,4096,4215,4337,4461,4586,4714,
									4845,4977,5111,5247,5386,5526,5668,5813,
									5959,6107,6256,6408,6561,6716,6872,7030,
									7189,7350,7512,7675,7840,8005,8172,8340,
									8508,8678,8848,9018,9190,9361,9533,9705,
									9878,10050,10222,10394,10566,10738,10908,
									11079,11248,11417,11585,11752,11917,12082,
									12244,12406,12565,12723,12879,13033,13185,
									13334,13482,13626,13769,13908,14045,14178,
									14309,14437,14561,14682,14799,14913,15024,
									15130,15233,15332,15427,15518,15604,15687,
									15765,15838,15908,15972,16032,16088,16139,
									16185,16227,16263,16295,16322,16344,16361,
									16374,16381,16384);
begin
	o_Data <= std_logic_vector(to_unsigned(values(to_integer(unsigned(i_Data))),g_bits));
end RTL;